module branch_control
(
  // current pc
  input branch,
  input check,

  output reg taken 
);

///////////////////////////////////////////////////////////////////////////////
// TODO : You need to do something!
//////////////////////////////////////////////////////////////////////////////
always @(*) begin
  taken = ({branch, check}==2'b11)? 1'b1:1'b0;
end
endmodule
